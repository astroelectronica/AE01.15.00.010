.title KiCad schematic
V1 /IN 0 AC 1
R1 0 /OUT {RHPF}
C1 /IN /OUT {CHPF}
.end
